library verilog;
use verilog.vl_types.all;
entity Golombtester is
end Golombtester;
